module test_verilog(
					input [17:0] SW,
					input CLOCK_50,
					output [17:0] LEDR,
					output [7:0] LEDG,
					output [6:0] HEX0,
					output [6:0] HEX1,
					output [6:0] HEX2,
					output [6:0] HEX3,
					output [6:0] HEX4,
					output [6:0] HEX5,
					output [6:0] HEX6,
					output [6:0] HEX7
					);


					%%PLACEHOLDER%%
	

endmodule
